library	IEEE;
use		IEEE.STD_LOGIC_1164		.all;
use		IEEE.STD_LOGIC_ARITH	.all;
use		IEEE.STD_LOGIC_UNSIGNED	.all;
use		IEEE.Numeric_STD		.all;



entity sync_generator is
	generic
	(
		-- this values depend on the input clq frequency and
		-- scan frequency. The following are HSYNC ones
		-- for the 25 MHz clk and 60 Hz scan frequency

		-- how many pixel clock cycles are spent on the display surface
		t_display			: integer := 640;
		-- how many pixel clock cycles we wait before dropping SYNC current
		t_fp				: integer := 16;
		-- how many pixel clock cycles we wait before starting drawing
		t_bp				: integer := 16;
		-- how many pixel clock cycles are needed for the magnetic field to lapse
		t_pw				: integer := 64;
		
		counter_width		: integer := 10
	);
	port
	(
		clock_i				: in	std_logic; -- main clock
		reset_i				: in	std_logic; -- main reset
		enable_i			: in	std_logic; -- enable -- pixel clock/row clock
		
		sync_o				: out	std_logic; -- output of HSYNC
		sig_cycle_o			: out	std_logic; -- row clock -- enable for vsync
		
		en_draw_o			: out	std_logic; -- enable drawing (on display surface)
		pixel_pos_o			: out	std_logic_vector(counter_width - 1 downto 0)
	);
end sync_generator;



architecture Behavioral of sync_generator is

	signal scancounter		: std_logic_vector(counter_width - 1 downto 0);
	signal scancounter_reset: std_logic;

	signal sig_cycle		: std_logic;

	signal sig_sync_off		: std_logic;
	signal sig_sync_on		: std_logic;
	signal sig_display_off	: std_logic;
	signal sig_display_on	: std_logic;

	signal sync_on			: std_logic;
	signal draw_on			: std_logic;

begin
	sig_cycle_o				<= sig_cycle;
	sig_cycle				<= sig_display_on;

	scancounter_reset		<= reset_i or sig_cycle;
	pixel_pos_o				<= scancounter;


	-- start of count is at beginning of display
	Inst_sync_counter:		entity work.counter
	GENERIC MAP				(width => counter_width)
	PORT MAP
	(
		clock_i				=> clock_i,
		reset_i				=> scancounter_reset,
		count_enable_i		=> enable_i,
		count_o				=> scancounter
	);


	-- signals when we fall off display
	Inst_comparator_off_display: entity work.comparator
	PORT MAP
	(
		a_i					=> scancounter,
		b_i					=> std_logic_vector(to_unsigned(t_display, counter_width)),
		eq_o				=> sig_display_off
	);

	-- signals when we have to turn off SYNC
	Inst_comparator_off_fp: entity work.comparator
	PORT MAP
	(
		a_i					=> scancounter,
		b_i					=> std_logic_vector(to_unsigned(t_display + t_fp, counter_width)),
		eq_o				=> sig_sync_off
	);

	-- signals when to turn SYNC back on
	Inst_comparator_off_pw: entity work.comparator
	PORT MAP
	(
		a_i					=> scancounter,
		b_i					=> std_logic_vector(to_unsigned(t_display + t_fp + t_pw, counter_width)),
		eq_o				=> sig_sync_on
	);

	-- signals when we have to reset the count and start over
	Inst_comparator_cycle: entity work.comparator
	PORT MAP
	(
		a_i					=> scancounter,
		b_i					=> std_logic_vector(to_unsigned(t_display + t_fp + t_pw + t_bp, counter_width)),
		eq_o				=> sig_display_on
	);

	
	process (sig_display_on, sig_display_off, draw_on)
	begin
		if sig_display_on = '1' then
			en_draw_o			<= '1';
		elsif draw_on = '1' and sig_display_off = '0' then
			en_draw_o			<= '1';
		else
			en_draw_o			<= '0';
		end if;
	end process;


	process (sig_sync_on, sig_sync_off, sync_on)
	begin
		if (sig_sync_on = '1' or sync_on = '1') and sig_sync_off = '0' then
			sync_o				<= '1';
		else
			sync_o				<= '0';
		end if;
	end process;


	Inst_flip_flop_jk_sync: entity work.flip_flop_jk
	PORT MAP
	(
		clock_i				=> clock_i,
		reset_i				=> reset_i,
		j_i					=> sig_sync_on,
		k_i					=> sig_sync_off,
		q_o					=> sync_on
	);
	
	
	Inst_flip_flop_jk_draw: entity work.flip_flop_jk
	PORT MAP
	(
		clock_i				=> clock_i,
		reset_i				=> reset_i,
		j_i					=> sig_display_on,
		k_i					=> sig_display_off,
		q_o					=> draw_on
	);

end Behavioral;
